CSbiased0_9V-10uAVoIo
* file: CSbiased0_9V-10uAVoIo
* Spice circuit file
.include CMOS18TT.lib
M1 2 1 0 0 C18nmos W=220n L=180n
VdsQ 2 3 0.9
IdsQ 0 3 10u
VgsQ 1 4 0.643709
Vi   4 0 0
Io   0 3 0
.dc Io -20u 20u 1u
.end
