"Voltage amplifier with VCVS controller"
* file: vAmpBlack.cir
* SLiCAP circuit file
V1 1 0 {V_s}
R1 1 2 {R_s}
R2 3 0 {R_ell} 
E1 3 0 2 4 {A_v}
R3 3 4 {R_a}
R4 4 0 {R_b}
.end
