cfbVampExtended
* file: cfbVampExtended.cir
* SLiCAP circuit file
V1 1 0 {V_s}
R1 1 2 {R_s}
O1 2 4 3 0 mycfb
R2 3 0 {R_ell}
R3 3 4 {R_a}
R4 4 0 {R_b}
* Model definition for the operational amplifier 'mycfb'
.model mycfb OC cp={C_i} gp={1/R_i} cpn={C_d} gpn={1/R_d} gm={g_m} 
+               zt={R_t/(1+s*tau)} zo={R_o/(1+s*tau)}
* parameter values for numeric simulation
.param C_i=5p R_i=1M g_m=20m R_t=1M R_o=2k tau=50u R_a=2k R_b=500 R_s=100
+             R_ell=500 V_s=1 C_d=2p R_d=10k
.end