* C:\Users\User\OneDrive\Documents\GitHub\SLiCAP_python\files\examples\Chapter5\SLiCAP\cir\shuntswitch_imp.asc
R1 N001 0 {R_L} noisetemp=0 noiseflow=0 dcvar=0
R3 source 0 {R_S} noisetemp=0 dcvar=0
I1 0 source I value=0 dc=0 dcvar=0 noise=0
I2 0 N001 I value=0 dc=0 dcvar=0 noise=0
C1 source P001 {Csb} vinit=0
C2 N001 P002 {Cdb} vinit=0
R2 P001 0 {Rb1}
R4 P002 0 {Rb2}
R5 N001 source {Rch}
C3 N001 source {Cch} vinit=0
.backanno
.end
