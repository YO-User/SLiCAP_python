"Root Locus 2nd order voltage amplifier"
* File: RLvAmp-2.cir
* SLiCAP netlist file
V1 1 0 {V_s}
R1 1 2 {R_s}
E1 3 0 2 4 {A_0/(1-s/p_1)/(1-s/p_2)}
E2 4 0 3 0 {A*(1-s/z_1)}
R2 3 0 {R_ell}
* For pole-zero analysis all parameters must have a numeric value
.param A_0 = 1M A = 10m
+ p_1 = {-2*pi} 
+ p_2 = {-2*pi*100} 
+ z_1 = {-2*pi*761.49}
+ R_ell = 1 R_s=1 V_s=1
.end
