RL1_L
* file: RL1_L.cir
V1 1 0 0
E1 2 0 1 2 {A_0*(1-s/2/pi/z_1)/(1-s/2/pi/p_1)}
.param A_0=100 p_1=-10 z_1=-100
.end