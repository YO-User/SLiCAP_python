"CS stage MOS small-signal model"
* Z:\mnt\DATA\Cursussen\Publish\Books\CSstage\SLiCAP\cir\CSstageModel.asc
R1 out 0 {R_L}
I1 0 N001 I value=0 dc=0 dcvar=0 noise=0
R2 N001 0 {R_s}
M1 out N001 0 0 myNMOS
.model myNMOS  M gm={g_m} cgs={c_gs} cgb={c_gb} cdg={c_dg} cdb={c_db} go={g_o}
.param R_s=10G R_L=10k
.backanno
.end
