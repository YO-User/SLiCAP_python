* C:\Users\User\OneDrive\Documents\GitHub\SLiCAP_python\files\examples\Chapter5\SLiCAP\cir\halfswitch_LKY.asc
R1 out2 0 {R_L} noisetemp=0 noiseflow=0 dcvar=0
R3 source 0 {R_S} noisetemp=0 dcvar=0
I1 0 source I value=0 dc=0 dcvar=0 noise=0
L2 N001 P001 {La} iinit=0
XU3 out2 0 in2 0 ABCD A={A2} B={B2} C={C2} D={D2}
I2 0 out2 I value=0 dc=0 dcvar=0 noise=0
XU1 out1 0 source 0 ABCD
L1 out1 0 {L1} iinit=0
L4 N003 N002 {Lb} iinit=0
C3 out1 P001 {ca} vinit=0
C1 out2 N002 {cb} vinit=0
R5 N001 in2 {ra} noisetemp=0 dcvar=0
R6 N003 0 {rb} noisetemp=0 dcvar=0
.model myNMOS  M gm={g_m} cgs={c_gs} cgb={c_gb} cdg={c_dg} cdb={c_db} go={g_o}
.param R_S=10G R_L=10k R_f=50 R_b=1.5k Z1=50 T1=10n Z2=50 T2=10n L=1n R7_comp=50 R8_comp=50
.model myNMOS2  M gm={g_mp} cgs={c_gsp} cgb={c_gbp} cdg={c_dgp} cdb={c_dbp} go={g_op}
.backanno
.end
