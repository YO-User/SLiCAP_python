* Sub circuit nNoise
* LTspice subcircuit for a noisy nullor for noise analysis
* Lowest frequency 100uHz
* For lower frequencies increase C1 and C2
* Nodes:       in+ in- out+ out- 
.subckt nNoise inP inN outP outN params: Sv=1n Si=1p flv=1k fli=10k
* Parameters:
* Sv:  input noise voltage density (noise-floor) in V/sqrt(Hz)
* flv: 1/f corner frequency of voltage noise
* Si:  input noise current density (noise-floor) in A/sqrt(Hz)
* fli: 1/f corner frequency of current noise
E1 outP 6 inP 5 1
E2 outP outN 6 outN 1
D1 1 3 DnoiseV
D2 3 outN DnoiseI
I1 outN 1 3.125u
C1 1 2 1
C2 3 4 1
Vi 2 3 0
Vv 4 outN 0
F1 inP inN Vi {Si*1e12}
H1 inN 5 Vv {Sv*1e12}
.model DnoiseV D kf={3.2e-19*flv} af=1
.model DnoiseI D kf={3.2e-19*fli} af=1
.ends nNoise
