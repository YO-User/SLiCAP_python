* C:\Users\User\OneDrive\Documents\GitHub\SLiCAP_python\files\examples\Chapter5\SLiCAP\cir\halfswitch_simp_A.asc
R1 out 0 {R_L} noisetemp=0 noiseflow=0 dcvar=0
M1 out N001 N002 N003 myNMOS
R3 source 0 {R_S} noisetemp=0 dcvar=0
I1 0 source I value=0 dc=0 dcvar=0 noise=0
R2 N003 0 {R_b}
R4 v1a N001 {R_b}
L2 out N002 {L} iinit=0
V1 v1a 0 V value=0 dc=0 dcvar=0 noise=0
XU1 N002 0 source 0 ABCD
L1 N002 0 {L1} iinit=0
I2 0 out I value=0 dc=0 dcvar=0 noise=0
.model myNMOS  M gm={g_m} cgs={c_gs} cgb={c_gb} cdg={c_dg} cdb={c_db} go={g_o}
.param R_S=10G R_L=10k R_f=50 R_b=1.5k Z1=50 T1=10n Z2=50 T2=10n L=1n R7_comp=50 R8_comp=50
.model myNMOS2  M gm={g_mp} cgs={c_gsp} cgb={c_gbp} cdg={c_dgp} cdb={c_dbp} go={g_op}
.backanno
.end
