"NA-2"
* file: NA-2.cir
* SLiCAP netlist for nodal analysis
I1 1 0 {I_s}
C1 0 1 {C_a}
R1 0 1 {R_a}
R2 0 2 {R_b}
C2 2 1 {C_b}
.param R_a=100k R_b=1k C_a=100p C_b=10n I_s=1
.end
