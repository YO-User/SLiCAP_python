R_3_0
* file: R_3_0.cir
V1 1 0 0
E1 2 0 1 2 {A_0/(20k*pi^2 + 200*pi*s + s^2)/s}
.param A_0 = 50
.end