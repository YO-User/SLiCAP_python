cfbVamp 
* file: cfbVamp.cir
* SLiCAP circuit file
V1 1 0 {V_s}
R1 1 2 {R_s}
R2 4 0 {R_ell}
R3 4 5 {R_a}
R4 5 0 {R_b}
G1 3 5 2 5 {g_m}
H1 4 0 0 3 H value={A_r}
.end
