myNPN_FT
* FILE: myNPN_FT.cir
* LTspice circuit file for plotting fT(Ic)
V1 4 1 3
V2 2 3 DC 0 AC 1
I1 0 4 {Ic}
C1 1 0 1
E1 2 0 1 0 1
Q1 4 3 0 myNPN
.model myNPN NPN
+ IS=0.5f BF=100 NF=1 IKF=100m ISE=10f NE=2 RB=10
+ TF=1n CJE=5p CJC=1p VJE=0.6 VJC=0.8 XTF=1 VTF=2 ITF=20m
.ac dec 50 1 1G
* LTspice syntax for plotting fT(Ic)
.step dec param Ic 100n 10m 10
.meas AC fT FIND Frequency WHEN dB(I(V1)/I(V2))=0 CROSS=1
* Run this netlist and press CTRL + L in the trace window
* This will bring up the output file (Spice error log) window
* In this window right-click "Plot .step'ed .meas data"
.end
