transimpedancePZcancel
* file: transimpedancePZcancel.cir
* SLiCAP circuit file
I1 0 1 0
C1 1 0 {C_s}
C2 1 0 {C_d}
C3 1 0 {C_c/2}
C4 3 0 {C_z}
R1 1 2 {R_f}
R2 2 0 {R_ell}
R3 1 3 {R_z}
E1 2 0 0 1 EZ value={A_0/(1+s/2/pi/16)} zo={R_o}
.param C_s=5p R_f=100k R_ell=2k C_d=8p C_c=7p A_0=1M 
+ R_o=55 C_z={1/R_z/2/pi/16} R_z=5.896k
.end
