* file: nullor.cir
* LTspice nullor subcircuit
.subckt nullor 3 4 1 2
E1 3 4 3 5 1
E2 5 4 1 2 1
.ends nullor