mosEKVplots
* SLiCAP netlist file
.include C18.lib
X1 d g s 0 CMOS18N W={W} L={L} ID={I_D}
.param I_D=1a W=220n L=180n
.end
