RL1_R
* file: RL1_R.cir
V1 1 0 0
E1 2 0 1 2 {A_0*(1-s/2/pi/z_1)/(1-s/2/pi/p_1)}
.param A_0=100 p_1=-100 z_1=-10
.end