VampNoise.cir
X1 2 3 out 0 N_noise si={S_i} sv={S_v}
R1 out 3 {R_b}
R2 3 0 {R_a}
I1 out 3 I noise={4*k*T/R_b}
I2 3 0 I noise={4*k*T/R_a}
R3 2 1 {R_s}
V1 1 0 V noise={4*k*T*R_s}
.end
