RL2_0
* file: RL2_0.cir
V1 1 0 0
E1 2 0 1 2 {A_0/(1-s/2/pi/p_1)/(1-s/2/pi/p_2)}
.param A_0=100 p_1=-10 p_2=-40
.end