* C:\Users\User\Documents\GitHub\SLiCAP_python\files\examples\Chapter5\SLiCAP\cir\CSstageModel4.asc
R1 out 0 {R_L} noisetemp=0 noiseflow=0 dcvar=0
M1 out N001 0 0 myNMOS
V1 N003 0 V value=0 dc=0 dcvar=0 noise=0
R3 N001 N003 {R_S} noisetemp=0 dcvar=0
M2 out N001 0 N002 myPMOS
R2 out N001 {R_f} noisetemp=0 dcvar=0
.model myNMOS  M gm={g_m} cgs={c_gs} cgb={c_gb} cdg={c_dg} cdb={c_db} go={g_o}
.param R_s=50 R_L=10k R_f=50
.model myPMOS  M gm={g_mp} cgs={c_gsp} cgb={c_gbp} cdg={c_dgp} cdb={c_dbp} go={g_op}
.backanno
.end
