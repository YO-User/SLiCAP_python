transimpedanceCompensatedSource
* file: transimpedanceCompensatedSource.cir
* SLiCAP circuit file
I1 0 1 0
C1 1 0 {C_s}
C2 3 0 {C_d}
C3 3 0 {C_c/2}
R1 3 2 {R_f}
R2 2 0 {R_ell}
R3 1 3 r value={R_phz}
E1 2 0 0 3 EZ value={A_0/(1+s*A_0/2/pi/G_B)} zo={R_o}
.param C_s=5p R_f=100k R_ell=2k C_d=8p C_c=7p A_0=1M R_o=55 G_B=16M R_phz=0
.end
